module diag

fn test_diag_ones_k_pos() {
	m := 7
	n := 4
	k := 5
	b := diag_ones(m, n, k)
	assert b == [0.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0,
		0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0]
	m_1 := 7
	n_1 := 4
	k_1 := 1
	b_1 := diag_ones(m_1, n_1, k_1)
	assert b_1 == [0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0,
		0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0]
	m_2 := 4
	n_2 := 7
	k_2 := 1
	b_2 := diag_ones(m_2, n_2, k_2)
	assert b_2 == [0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0,
		0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0]
	m_3 := 4
	n_3 := 4
	k_3 := 0
	b_3 := diag_ones(m_3, n_3, k_3)
	assert b_3 == [1.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 1.0]
}

fn test_diag_ones_k_neg() {
	m := 7
	n := 5
	k := -1
	b := diag_ones(m, n, k)
	assert b == [0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 1.0,
		0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0,
		0.0]
	m_1 := 4
	n_1 := 7
	k_1 := -1
	b_1 := diag_ones(m_1, n_1, k_1)
	assert b_1 == [0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0,
		0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0]
	m_2 := 4
	n_2 := 4
	k_2 := -1
	b_2 := diag_ones(m_2, n_2, k_2)
	assert b_2 == [0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0]
}

fn test_diag_arb_k_pos() {
	m := 7
	n := 4
	k := 5
	val := [1.0, 2.0]
	b := diag_arb(m, n, k, val)
	assert b == [0.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 2.0, 0.0, 0.0,
		0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0]
	m_1 := 7
	n_1 := 4
	k_1 := 1
	val_1 := [1.0, 2.0, 3.0, 4.0]
	b_1 := diag_arb(m_1, n_1, k_1, val_1)
	assert b_1 == [0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 2.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0,
		0.0, 3.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 4.0, 0.0, 0.0]
	m_2 := 4
	n_2 := 7
	k_2 := 1
	val_2 := [1.0, 2.0, 3.0]
	b_2 := diag_arb(m_2, n_2, k_2, val_2)
	assert b_2 == [0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 2.0, 0.0, 0.0, 0.0, 0.0, 3.0, 0.0, 0.0, 0.0, 0.0,
		0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0]
	m_3 := 4
	n_3 := 4
	k_3 := 0
	val_3 := [1.0, 2.0, 3.0, 4.0]
	b_3 := diag_arb(m_3, n_3, k_3, val_3)
	assert b_3 == [1.0, 0.0, 0.0, 0.0, 0.0, 2.0, 0.0, 0.0, 0.0, 0.0, 3.0, 0.0, 0.0, 0.0, 0.0, 4.0]
}

fn test_diag_arb_k_neg() {
	m := 7
	n := 5
	k := -1
	val := [1.0, 2.0, 3.0, 4.0]
	b := diag_arb(m, n, k, val)
	assert b == [0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 2.0,
		0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 3.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 4.0, 0.0, 0.0,
		0.0]
	m_1 := 4
	n_1 := 7
	k_1 := -1
	val_1 := [1.0, 2.0, 3.0, 4.0]
	b_1 := diag_arb(m_1, n_1, k_1, val_1)
	assert b_1 == [0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 2.0, 0.0, 0.0, 0.0, 0.0, 3.0, 0.0,
		0.0, 0.0, 0.0, 4.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0]
	m_2 := 4
	n_2 := 4
	k_2 := -1
	val_2 := [1.0, 2.0, 3.0]
	b_2 := diag_arb(m_2, n_2, k_2, val_2)
	assert b_2 == [0.0, 0.0, 0.0, 0.0, 1.0, 0.0, 0.0, 0.0, 0.0, 2.0, 0.0, 0.0, 0.0, 0.0, 3.0, 0.0]
}

